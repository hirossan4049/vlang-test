module testmodule


pub fn test() {
	println("hey, Python! I'm V-lang!")
}
